.title KiCad schematic
.include "C:/AE/LT1762/_models/C3216X5R2A105K160AA_s.mod"
.include "C:/AE/LT1762/_models/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/LT1762/_models/CGA5L3X5R1H106K160AB_s.mod"
.include "C:/AE/LT1762/_models/LT1762.lib"
R2 /VOUT /ADJ {RADJU}
XU3 /BYP /VOUT CEU4J2X7R2A103K125AE_s
R3 /ADJ 0 {RADJB}
I1 /VOUT 0 {ILOAD}
XU4 /VOUT 0 CGA5L3X5R1H106K160AB_s
XU1 /VIN 0 C3216X5R2A105K160AA_s
V1 /VIN 0 {VSOURCE}
XU2 /VOUT /ADJ /BYP 0 /VIN /VIN LT1762
.end
